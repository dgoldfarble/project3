module RF	(	// inputs
				//outputs
			);
			
	
	output reg      [31: 0] Reg [0:31];
